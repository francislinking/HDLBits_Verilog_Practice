module top_module (
	input clk,
	input resetn,
	input in,
	output out
);

	reg [3:0] sr;
	
	// Create a shift register named sr. It shifts in "in".
	always @(posedge clk) begin
		if (~resetn)		// Synchronous active-low reset
			sr <= 0;
		else 
			sr <= {sr[2:0], in};
	end
	
	assign out = sr[3];		// Output the final bit (sr[3])


    // my solution
    // reg [2:0] Q;
    // always @ (posedge clk) begin
    //     if (~resetn)
    //     	{out,Q}<=4'h0;
    //     else
    //     	{out,Q}<={Q,in};   
    // end
    
endmodule
