module top_module (
    input d, 
    input ena,
    output q);
	
    always @(ena) begin
        q = ena? d : q;
    end
endmodule
