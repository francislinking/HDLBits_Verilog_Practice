module top_module(
	input clk,
	input load,
	input [511:0] data,
	output reg [511:0] q);
	
	always @(posedge clk) begin
		if (load)
			q <= data;	// Load the DFFs with a value.
		else begin
			// At each clock, the DFF storing each bit position becomes the XOR of its left neighbour
			// and its right neighbour. Since the operation is the same for every
			// bit position, it can be written as a single operation on vectors.
			// The shifts are accomplished using part select and concatenation operators.
			
			//     left           right
			//  neighbour       neighbour
			q <= q[511:1] ^ {q[510:0], 1'b0} ;
		end
	end

    // my solution
    // wire [511:0] L,R;
    // assign L = {1'b0,q[511:1]};
    // assign R = {q[510:0],1'b0};
    
    // always @(posedge clk) begin
    //     if (load)
    //         q<=data;
    //     else begin
    //         q<=L^R;
    //     end
    // end


endmodule
